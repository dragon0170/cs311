module ImmediateGenerator(input [31:0] part_of_inst, output [31:0] imm_gen_out);
  
endmodule